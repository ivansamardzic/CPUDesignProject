module shr_32_bit(input wire [31:0] in, [31:0] shift, output wire[31:0] out);

assign out = in >> shift; 

endmodule
